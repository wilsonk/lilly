module buffer

import arrays

pub struct GapBuffer {
mut:
	buffer       []rune
	pre_gap_len  int
	post_gap_len int
}

const c_gapsize = 50

pub fn new_gap_buffer(size int) &GapBuffer {
	mut len := size - c_gapsize
	if len < c_gapsize { len = c_gapsize }
	return &GapBuffer{ buffer: []rune{ len: len, cap: len } }
}

pub fn (mut gap_buffer GapBuffer) set_string(s string) {
	gap_buffer.buffer = s.runes()
	gap_buffer.pre_gap_len = 0
	gap_buffer.post_gap_len = gap_buffer.buffer.len
	gap_buffer.move_cursor_left()
}

pub fn (mut gap_buffer GapBuffer) get_string() string {
	mut text := []rune{}
	text << gap_buffer.buffer[..gap_buffer.pre_gap_len]
	text << gap_buffer.buffer[gap_buffer.post_gap_start()..]
	return text.string()
}

/*
// moveGap moves the gap to the specified position.
func (gb *GapBuffer) moveGap(pos int) {
	gapStart := gb.gapPos
	gapEnd := gb.gapPos + gb.gapLen
	copy(gb.buf[pos+gb.gapLen:], gb.buf[gapEnd:])
	copy(gb.buf[pos:], gb.buf[gapStart:gapEnd])
	gb.gapPos = pos
}
*/

pub fn (mut gap_buffer GapBuffer) move_cursor_left() bool {
	if gap_buffer.pre_gap_len == 0 { return false }
	gap_buffer.buffer[gap_buffer.post_gap_start() - 1] = gap_buffer.buffer[gap_buffer.pre_gap_len - 1]
	gap_buffer.pre_gap_len -= 1
	gap_buffer.post_gap_len += 1
	return true
}

pub fn (mut gap_buffer GapBuffer) move_cursor_right() bool {
	if gap_buffer.post_gap_len == 0 { return false }
	gap_buffer.buffer[gap_buffer.pre_gap_len] = gap_buffer.buffer[gap_buffer.post_gap_start()]
	gap_buffer.pre_gap_len += 1
	gap_buffer.post_gap_len -= 1
	return true
}

pub fn (mut gap_buffer GapBuffer) insert(c rune) {
	if gap_buffer.gap_len() == 0 {
		gap_buffer.grow_gap()
	}
	gap_buffer.buffer[gap_buffer.gap_start()] = c
	gap_buffer.pre_gap_len += 1
}

pub fn (mut gap_buffer GapBuffer) delete() bool {
	if gap_buffer.post_gap_len == 0 { return false }
	gap_buffer.post_gap_len -= 1
	return true
}

pub fn (mut gap_buffer GapBuffer) backspace() bool {
	if gap_buffer.pre_gap_len == 0 { return false }
	gap_buffer.pre_gap_len -= 1
	return true
}

fn (mut gap_buffer GapBuffer) get_line_str(line_num int) !string {
	if line_num < 0 { return error("invalid line index ${line_num} < 0") }
	newline_locations := gap_buffer.locate_newlines()
	if line_num > newline_locations.len { return error("invalid line index ${line_num} > ${newline_locations.len}") }

	// FIX(tauraamui): don't really want to do this, it's probably creating a copy, look into direct access more
	mut document := gap_buffer.buffer[..gap_buffer.pre_gap_len]
	document << gap_buffer.buffer[gap_buffer.post_gap_start()..]

	if newline_locations.len == 0 {
		if line_num == 0 { return document.string() }
		return error("invalid line index ${line_num > 0}")
	}

	// if want to retrieve line 0/1
	if line_num == 0 {
		return document[..newline_locations[0]].string()
	}

	// if want to retrieve last line
	if line_num == newline_locations.len {
		return document[newline_locations[line_num - 1] + 1..].string()
	}

	return document[newline_locations[line_num - 1] + 1..newline_locations[line_num]].string()
}

fn (mut gap_buffer GapBuffer) get_lines_str(from int, to int) []string {
	mut lines := []string{}
	for i := from; i <= to; i++ {
		lines << gap_buffer.get_line_str(i) or { continue }
	}
	return lines
}

fn (mut gap_buffer GapBuffer) locate_newlines() []int {
	mut found := []int{}
	for i, r in gap_buffer.buffer[..gap_buffer.pre_gap_len] { if r == `\n` { found << i } }
	for i, r in gap_buffer.buffer[gap_buffer.post_gap_start()..] { if r == `\n` { found << i + gap_buffer.gap_len() } }
	return found
}

// TODO(tauraamui) -> use this at some point
fn (mut gap_buffer GapBuffer) locate_newlines_2() ([]int, []int) {
	mut pre_gap_found := []int{}
	mut post_gap_found := []int{}

	for i, r in gap_buffer.buffer[..gap_buffer.pre_gap_len] { if r == `\n` { pre_gap_found << i } }
	for i, r in gap_buffer.buffer[gap_buffer.post_gap_start()..] { if r == `\n` { post_gap_found << i + gap_buffer.gap_len() } }

	return pre_gap_found, post_gap_found
}

fn (mut gap_buffer GapBuffer) gap_start() int {
	return gap_buffer.pre_gap_len
}

fn (mut gap_buffer GapBuffer) gap_len() int {
	return gap_buffer.post_gap_start() - gap_buffer.pre_gap_len
}

fn (mut gap_buffer GapBuffer) post_gap_start() int {
	return gap_buffer.buffer.len - gap_buffer.post_gap_len
}

fn (mut gap_buffer GapBuffer) grow_gap() {
	mut new_buffer := []rune{ len: gap_buffer.buffer.len * 2, cap: gap_buffer.buffer.len * 2 }
	arrays.copy(mut &new_buffer, gap_buffer.buffer[..gap_buffer.pre_gap_len])
	new_buffer.insert(gap_buffer.post_gap_start(), gap_buffer.buffer[gap_buffer.post_gap_start()..])
	gap_buffer.buffer = new_buffer
}

