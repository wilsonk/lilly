module piece_tree

fn test_alloc() {
	p := Piece{}
	assert p == Piece{}
}
