module piece_tree

struct UndoRedoEntry {
}
