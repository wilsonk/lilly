module piece_tree

fn test_alloc() {
	r := new_tree()
}
